library ieee;
use ieee.std_logic_1164.all;

--entity extender_8to16 is
    --generic(
        --operand_width : integer:=16
        --);
    --port (
        --A: in std_logic_vector(7 downto 0);
        --B: out std_logic_vector(operand_width-1 downto 0)
    --) ;
--end extender_8to16;


entity extender_9to16 is
    generic(
        operand_width : integer:=16
        );
    port (
        A: in std_logic_vector(8 downto 0);
		  sel: in std_logic;
        B: out std_logic_vector(operand_width-1 downto 0)
    ) ;
end extender_9to16;


entity extender_6to16 is
    generic(
        operand_width : integer:=16
        );
    port (
        A: in std_logic_vector(5 downto 0);
        B: out std_logic_vector(operand_width-1 downto 0)
    ) ;
end extender_6to16;

--architecture a1 of extender_8to16 is
    
--begin
--shift8to16 : process( A, B )
--begin
			--B <= "00000000"&A;
		
--end process ; -- shift8to16
--end a1 ; -- a1


architecture a2 of extender_9to16 is
    
begin
shift9to16 : process( A, B, sel )
begin
		if (sel = "0") then 
			B <= "0000000"&A;						--Zero at MSB
		else 
			B <= A&"0000000";						--Zero at LSB
		end if;
		
end process ; -- shift9to16

signal pc, RF_d1, RF_d2, RF_d3, ls_out, seB, t2, t1, aluA, aluB, aluC: std_logic_vector(15 downto 0);
begin
ext1 : process( A,B,sel )
begin
if (controlword_SE2="01") then
    A <= IR(8 downto 0);
    B <= RF_d3;
    sel <= "1";
elsif (controlword_SE2="10") then
    A <= IR(8 downto 0);
    B <= aluB;
    sel <= "0";
end a2 ; -- a1


architecture a3 of extender_6to16 is
    
begin
shift6to16 : process( A, B )
begin
			B <= "0000000000"&A;
		
end process ; -- shift6to16

signal pc, RF_d1, RF_d2, ls_out, seB, t2, t1: std_logic_vector(15 downto 0);
begin
ext2 : process( A,B )
begin
if (controlword_SE1="01") then
    A <= IR(5 downto 0);
    B <= aluB;
if (controlword_SE1="10") then
    A <= IR(5 downto 0);
    B <= aluA;
end a3 ; -- a1
